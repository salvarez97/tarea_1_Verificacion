//compuerta and 2 entradas
module and2(
    input a,
    input b,
    output y
);

assign y = a & b;
endmodule